----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Sean Conway
-- 
-- Create Date: 09.10.2023 08:44:27
-- Design Name: 
-- Module Name: RF_Mux32_32Bit_22335824 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity RF_Mux32_32Bit_22335824 is
    port ( I0, I1, I2, I3 : in std_logic_vector (31 downto 0);
           I4, I5, I6, I7 : in std_logic_vector (31 downto 0);
           I8, I9, I10, I11 : in std_logic_vector (31 downto 0);
           I12, I13, I14, I15 : in std_logic_vector (31 downto 0);
           I16, I17, I18, I19 : in std_logic_vector (31 downto 0);
           I20, I21, I22, I23 : in std_logic_vector (31 downto 0);
           I24, I25, I26, I27 : in std_logic_vector (31 downto 0);
           I28, I29, I30, I31 : in std_logic_vector (31 downto 0);
           S : in std_logic_vector (4 downto 0);
           Y : out std_logic_vector (31 downto 0));
end RF_Mux32_32Bit_22335824;

architecture Behavioral of RF_Mux32_32Bit_22335824 is

        component RF_Mux32_1Bit_22335824
        port (I: in std_logic_vector (31 downto 0);
           S: in std_logic_vector (4 downto 0);
           Y: out std_logic
           );
        end component;
           
        constant AND_gate_delay : Time := 5ns;      -- least significant digit 5 = 4 + 1
        constant NAND_gate_delay : Time := 3ns;     -- next more significant digit 3 = 2 + 1
        constant OR_gate_delay : Time := 9ns;       -- next more significant digit 9 = 8 + 1
        constant NOR_gate_delay : Time := 6ns;      -- next more significant digit 6 = 5 + 1
        constant XOR_gate_delay : Time := 4ns;      -- next more significant digit 4 = 3 + 1
        constant XNOR_gate_delay : Time := 4ns;     -- next more significant digit 4 = 3 + 1
        constant NOT_gate_delay : Time := 3ns;      -- next more significant digit 3 = 2 + 1

begin

    bit0: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(0), I(1) => I1(0), I(2) => I2(0), I(3) => I3(0),
    I(4) => I4(0), I(5) => I5(0), I(6) => I6(0), I(7) => I7(0),
    I(8) => I8(0), I(9) => I9(0), I(10) => I10(0), I(11) => I11(0),
    I(12) => I12(0), I(13) => I13(0), I(14) => I14(0), I(15) => I15(0),
    I(16) => I16(0), I(17) => I17(0), I(18) => I18(0), I(19) => I19(0),
    I(20) => I20(0), I(21) => I21(0), I(22) => I22(0), I(23) => I23(0),
    I(24) => I24(0), I(25) => I25(0), I(26) => I26(0), I(27) => I27(0),
    I(28) => I28(0), I(29) => I29(0), I(30) => I30(0), I(31) => I31(0),
    S => S, Y => Y(0));
    
    bit1: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(1), I(1) => I1(1), I(2) => I2(1), I(3) => I3(1),
    I(4) => I4(1), I(5) => I5(1), I(6) => I6(1), I(7) => I7(1),
    I(8) => I8(1), I(9) => I9(1), I(10) => I10(1), I(11) => I11(1),
    I(12) => I12(1), I(13) => I13(1), I(14) => I14(1), I(15) => I15(1),
    I(16) => I16(1), I(17) => I17(1), I(18) => I18(1), I(19) => I19(1),
    I(20) => I20(1), I(21) => I21(1), I(22) => I22(1), I(23) => I23(1),
    I(24) => I24(1), I(25) => I25(1), I(26) => I26(1), I(27) => I27(1),
    I(28) => I28(1), I(29) => I29(1), I(30) => I30(1), I(31) => I31(1),
    S => S, Y => Y(1));
    
    bit2: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(2), I(1) => I1(2), I(2) => I2(2), I(3) => I3(2),
    I(4) => I4(2), I(5) => I5(2), I(6) => I6(2), I(7) => I7(2),
    I(8) => I8(2), I(9) => I9(2), I(10) => I10(2), I(11) => I11(2),
    I(12) => I12(2), I(13) => I13(2), I(14) => I14(2), I(15) => I15(2),
    I(16) => I16(2), I(17) => I17(2), I(18) => I18(2), I(19) => I19(2),
    I(20) => I20(2), I(21) => I21(2), I(22) => I22(2), I(23) => I23(2),
    I(24) => I24(2), I(25) => I25(2), I(26) => I26(2), I(27) => I27(2),
    I(28) => I28(2), I(29) => I29(2), I(30) => I30(2), I(31) => I31(2),
    S => S, Y => Y(2));
    
    bit3: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(3), I(1) => I1(3), I(2) => I2(3), I(3) => I3(3),
    I(4) => I4(3), I(5) => I5(3), I(6) => I6(3), I(7) => I7(3),
    I(8) => I8(3), I(9) => I9(3), I(10) => I10(3), I(11) => I11(3),
    I(12) => I12(3), I(13) => I13(3), I(14) => I14(3), I(15) => I15(3),
    I(16) => I16(3), I(17) => I17(3), I(18) => I18(3), I(19) => I19(3),
    I(20) => I20(3), I(21) => I21(3), I(22) => I22(3), I(23) => I23(3),
    I(24) => I24(3), I(25) => I25(3), I(26) => I26(3), I(27) => I27(3),
    I(28) => I28(3), I(29) => I29(3), I(30) => I30(3), I(31) => I31(3),
    S => S, Y => Y(3));
    
    bit4: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(4), I(1) => I1(4), I(2) => I2(4), I(3) => I3(4),
    I(4) => I4(4), I(5) => I5(4), I(6) => I6(4), I(7) => I7(4),
    I(8) => I8(4), I(9) => I9(4), I(10) => I10(4), I(11) => I11(4),
    I(12) => I12(4), I(13) => I13(4), I(14) => I14(4), I(15) => I15(4),
    I(16) => I16(4), I(17) => I17(4), I(18) => I18(4), I(19) => I19(4),
    I(20) => I20(4), I(21) => I21(4), I(22) => I22(4), I(23) => I23(4),
    I(24) => I24(4), I(25) => I25(4), I(26) => I26(4), I(27) => I27(4),
    I(28) => I28(4), I(29) => I29(4), I(30) => I30(4), I(31) => I31(4),
    S => S, Y => Y(4));
    
    bit5: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(5), I(1) => I1(5), I(2) => I2(5), I(3) => I3(5),
    I(4) => I4(5), I(5) => I5(5), I(6) => I6(5), I(7) => I7(5),
    I(8) => I8(5), I(9) => I9(5), I(10) => I10(5), I(11) => I11(5),
    I(12) => I12(5), I(13) => I13(5), I(14) => I14(5), I(15) => I15(5),
    I(16) => I16(5), I(17) => I17(5), I(18) => I18(5), I(19) => I19(5),
    I(20) => I20(5), I(21) => I21(5), I(22) => I22(5), I(23) => I23(5),
    I(24) => I24(5), I(25) => I25(5), I(26) => I26(5), I(27) => I27(5),
    I(28) => I28(5), I(29) => I29(5), I(30) => I30(5), I(31) => I31(5),
    S => S, Y => Y(5));
    
    bit6: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(6), I(1) => I1(6), I(2) => I2(6), I(3) => I3(6),
    I(4) => I4(6), I(5) => I5(6), I(6) => I6(6), I(7) => I7(6),
    I(8) => I8(6), I(9) => I9(6), I(10) => I10(6), I(11) => I11(6),
    I(12) => I12(6), I(13) => I13(6), I(14) => I14(6), I(15) => I15(6),
    I(16) => I16(6), I(17) => I17(6), I(18) => I18(6), I(19) => I19(6),
    I(20) => I20(6), I(21) => I21(6), I(22) => I22(6), I(23) => I23(6),
    I(24) => I24(6), I(25) => I25(6), I(26) => I26(6), I(27) => I27(6),
    I(28) => I28(6), I(29) => I29(6), I(30) => I30(6), I(31) => I31(6),
    S => S, Y => Y(6));
    
    bit7: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(7), I(1) => I1(7), I(2) => I2(7), I(3) => I3(7),
    I(4) => I4(7), I(5) => I5(7), I(6) => I6(7), I(7) => I7(7),
    I(8) => I8(7), I(9) => I9(7), I(10) => I10(7), I(11) => I11(7),
    I(12) => I12(7), I(13) => I13(7), I(14) => I14(7), I(15) => I15(7),
    I(16) => I16(7), I(17) => I17(7), I(18) => I18(7), I(19) => I19(7),
    I(20) => I20(7), I(21) => I21(7), I(22) => I22(7), I(23) => I23(7),
    I(24) => I24(7), I(25) => I25(7), I(26) => I26(7), I(27) => I27(7),
    I(28) => I28(7), I(29) => I29(7), I(30) => I30(7), I(31) => I31(7),
    S => S, Y => Y(7));
    
    bit8: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(8), I(1) => I1(8), I(2) => I2(8), I(3) => I3(8),
    I(4) => I4(8), I(5) => I5(8), I(6) => I6(8), I(7) => I7(8),
    I(8) => I8(8), I(9) => I9(8), I(10) => I10(8), I(11) => I11(8),
    I(12) => I12(8), I(13) => I13(8), I(14) => I14(8), I(15) => I15(8),
    I(16) => I16(8), I(17) => I17(8), I(18) => I18(8), I(19) => I19(8),
    I(20) => I20(8), I(21) => I21(8), I(22) => I22(8), I(23) => I23(8),
    I(24) => I24(8), I(25) => I25(8), I(26) => I26(8), I(27) => I27(8),
    I(28) => I28(8), I(29) => I29(8), I(30) => I30(8), I(31) => I31(8),
    S => S, Y => Y(8));
    
    bit9: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(9), I(1) => I1(9), I(2) => I2(9), I(3) => I3(9),
    I(4) => I4(9), I(5) => I5(9), I(6) => I6(9), I(7) => I7(9),
    I(8) => I8(9), I(9) => I9(9), I(10) => I10(9), I(11) => I11(9),
    I(12) => I12(9), I(13) => I13(9), I(14) => I14(9), I(15) => I15(9),
    I(16) => I16(9), I(17) => I17(9), I(18) => I18(9), I(19) => I19(9),
    I(20) => I20(9), I(21) => I21(9), I(22) => I22(9), I(23) => I23(9),
    I(24) => I24(9), I(25) => I25(9), I(26) => I26(9), I(27) => I27(9),
    I(28) => I28(9), I(29) => I29(9), I(30) => I30(9), I(31) => I31(9),
    S => S, Y => Y(9));
    
    bit10: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(10), I(1) => I1(10), I(2) => I2(10), I(3) => I3(10),
    I(4) => I4(10), I(5) => I5(10), I(6) => I6(10), I(7) => I7(10),
    I(8) => I8(10), I(9) => I9(10), I(10) => I10(10), I(11) => I11(10),
    I(12) => I12(10), I(13) => I13(10), I(14) => I14(10), I(15) => I15(10),
    I(16) => I16(10), I(17) => I17(10), I(18) => I18(10), I(19) => I19(10),
    I(20) => I20(10), I(21) => I21(10), I(22) => I22(10), I(23) => I23(10),
    I(24) => I24(10), I(25) => I25(10), I(26) => I26(10), I(27) => I27(10),
    I(28) => I28(10), I(29) => I29(10), I(30) => I30(10), I(31) => I31(10),
    S => S, Y => Y(10));
    
    bit11: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(11), I(1) => I1(11), I(2) => I2(11), I(3) => I3(11),
    I(4) => I4(11), I(5) => I5(11), I(6) => I6(11), I(7) => I7(11),
    I(8) => I8(11), I(9) => I9(11), I(10) => I10(11), I(11) => I11(11),
    I(12) => I12(11), I(13) => I13(11), I(14) => I14(11), I(15) => I15(11),
    I(16) => I16(11), I(17) => I17(11), I(18) => I18(11), I(19) => I19(11),
    I(20) => I20(11), I(21) => I21(11), I(22) => I22(11), I(23) => I23(11),
    I(24) => I24(11), I(25) => I25(11), I(26) => I26(11), I(27) => I27(11),
    I(28) => I28(11), I(29) => I29(11), I(30) => I30(11), I(31) => I31(11),
    S => S, Y => Y(11));
    
    bit12: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(12), I(1) => I1(12), I(2) => I2(12), I(3) => I3(12),
    I(4) => I4(12), I(5) => I5(12), I(6) => I6(12), I(7) => I7(12),
    I(8) => I8(12), I(9) => I9(12), I(10) => I10(12), I(11) => I11(12),
    I(12) => I12(12), I(13) => I13(12), I(14) => I14(12), I(15) => I15(12),
    I(16) => I16(12), I(17) => I17(12), I(18) => I18(12), I(19) => I19(12),
    I(20) => I20(12), I(21) => I21(12), I(22) => I22(12), I(23) => I23(12),
    I(24) => I24(12), I(25) => I25(12), I(26) => I26(12), I(27) => I27(12),
    I(28) => I28(12), I(29) => I29(12), I(30) => I30(12), I(31) => I31(12),
    S => S, Y => Y(12));
    
    bit13: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(13), I(1) => I1(13), I(2) => I2(13), I(3) => I3(13),
    I(4) => I4(13), I(5) => I5(13), I(6) => I6(13), I(7) => I7(13),
    I(8) => I8(13), I(9) => I9(13), I(10) => I10(13), I(11) => I11(13),
    I(12) => I12(13), I(13) => I13(13), I(14) => I14(13), I(15) => I15(13),
    I(16) => I16(13), I(17) => I17(13), I(18) => I18(13), I(19) => I19(13),
    I(20) => I20(13), I(21) => I21(13), I(22) => I22(13), I(23) => I23(13),
    I(24) => I24(13), I(25) => I25(13), I(26) => I26(13), I(27) => I27(13),
    I(28) => I28(13), I(29) => I29(13), I(30) => I30(13), I(31) => I31(13),
    S => S, Y => Y(13));
    
    bit14: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(14), I(1) => I1(14), I(2) => I2(14), I(3) => I3(14),
    I(4) => I4(14), I(5) => I5(14), I(6) => I6(14), I(7) => I7(14),
    I(8) => I8(14), I(9) => I9(14), I(10) => I10(14), I(11) => I11(14),
    I(12) => I12(14), I(13) => I13(14), I(14) => I14(14), I(15) => I15(14),
    I(16) => I16(14), I(17) => I17(14), I(18) => I18(14), I(19) => I19(14),
    I(20) => I20(14), I(21) => I21(14), I(22) => I22(14), I(23) => I23(14),
    I(24) => I24(14), I(25) => I25(14), I(26) => I26(14), I(27) => I27(14),
    I(28) => I28(14), I(29) => I29(14), I(30) => I30(14), I(31) => I31(14),
    S => S, Y => Y(14));
    
    bit15: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(15), I(1) => I1(15), I(2) => I2(15), I(3) => I3(15),
    I(4) => I4(15), I(5) => I5(15), I(6) => I6(15), I(7) => I7(15),
    I(8) => I8(15), I(9) => I9(15), I(10) => I10(15), I(11) => I11(15),
    I(12) => I12(15), I(13) => I13(15), I(14) => I14(15), I(15) => I15(15),
    I(16) => I16(15), I(17) => I17(15), I(18) => I18(15), I(19) => I19(15),
    I(20) => I20(15), I(21) => I21(15), I(22) => I22(15), I(23) => I23(15),
    I(24) => I24(15), I(25) => I25(15), I(26) => I26(15), I(27) => I27(15),
    I(28) => I28(15), I(29) => I29(15), I(30) => I30(15), I(31) => I31(15),
    S => S, Y => Y(15));
    
    bit16: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(16), I(1) => I1(16), I(2) => I2(16), I(3) => I3(16),
    I(4) => I4(16), I(5) => I5(16), I(6) => I6(16), I(7) => I7(16),
    I(8) => I8(16), I(9) => I9(16), I(10) => I10(16), I(11) => I11(16),
    I(12) => I12(16), I(13) => I13(16), I(14) => I14(16), I(15) => I15(16),
    I(16) => I16(16), I(17) => I17(16), I(18) => I18(16), I(19) => I19(16),
    I(20) => I20(16), I(21) => I21(16), I(22) => I22(16), I(23) => I23(16),
    I(24) => I24(16), I(25) => I25(16), I(26) => I26(16), I(27) => I27(16),
    I(28) => I28(16), I(29) => I29(16), I(30) => I30(16), I(31) => I31(16),
    S => S, Y => Y(16));
    
    bit17: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(17), I(1) => I1(17), I(2) => I2(17), I(3) => I3(17),
    I(4) => I4(17), I(5) => I5(17), I(6) => I6(17), I(7) => I7(17),
    I(8) => I8(17), I(9) => I9(17), I(10) => I10(17), I(11) => I11(17),
    I(12) => I12(17), I(13) => I13(17), I(14) => I14(17), I(15) => I15(17),
    I(16) => I16(17), I(17) => I17(17), I(18) => I18(17), I(19) => I19(17),
    I(20) => I20(17), I(21) => I21(17), I(22) => I22(17), I(23) => I23(17),
    I(24) => I24(17), I(25) => I25(17), I(26) => I26(17), I(27) => I27(17),
    I(28) => I28(17), I(29) => I29(17), I(30) => I30(17), I(31) => I31(17),
    S => S, Y => Y(17));
    
    bit18: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(18), I(1) => I1(18), I(2) => I2(18), I(3) => I3(18),
    I(4) => I4(18), I(5) => I5(18), I(6) => I6(18), I(7) => I7(18),
    I(8) => I8(18), I(9) => I9(18), I(10) => I10(18), I(11) => I11(18),
    I(12) => I12(18), I(13) => I13(18), I(14) => I14(18), I(15) => I15(18),
    I(16) => I16(18), I(17) => I17(18), I(18) => I18(18), I(19) => I19(18),
    I(20) => I20(18), I(21) => I21(18), I(22) => I22(18), I(23) => I23(18),
    I(24) => I24(18), I(25) => I25(18), I(26) => I26(18), I(27) => I27(18),
    I(28) => I28(18), I(29) => I29(18), I(30) => I30(18), I(31) => I31(18),
    S => S, Y => Y(18));
    
    bit19: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(19), I(1) => I1(19), I(2) => I2(19), I(3) => I3(19),
    I(4) => I4(19), I(5) => I5(19), I(6) => I6(19), I(7) => I7(19),
    I(8) => I8(19), I(9) => I9(19), I(10) => I10(19), I(11) => I11(19),
    I(12) => I12(19), I(13) => I13(19), I(14) => I14(19), I(15) => I15(19),
    I(16) => I16(19), I(17) => I17(19), I(18) => I18(19), I(19) => I19(19),
    I(20) => I20(19), I(21) => I21(19), I(22) => I22(19), I(23) => I23(19),
    I(24) => I24(19), I(25) => I25(19), I(26) => I26(19), I(27) => I27(19),
    I(28) => I28(19), I(29) => I29(19), I(30) => I30(19), I(31) => I31(19),
    S => S, Y => Y(19));
    
    bit20: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(20), I(1) => I1(20), I(2) => I2(20), I(3) => I3(20),
    I(4) => I4(20), I(5) => I5(20), I(6) => I6(20), I(7) => I7(20),
    I(8) => I8(20), I(9) => I9(20), I(10) => I10(20), I(11) => I11(20),
    I(12) => I12(20), I(13) => I13(20), I(14) => I14(20), I(15) => I15(20),
    I(16) => I16(20), I(17) => I17(20), I(18) => I18(20), I(19) => I19(20),
    I(20) => I20(20), I(21) => I21(20), I(22) => I22(20), I(23) => I23(20),
    I(24) => I24(20), I(25) => I25(20), I(26) => I26(20), I(27) => I27(20),
    I(28) => I28(20), I(29) => I29(20), I(30) => I30(20), I(31) => I31(20),
    S => S, Y => Y(20));
    
    bit21: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(21), I(1) => I1(21), I(2) => I2(21), I(3) => I3(21),
    I(4) => I4(21), I(5) => I5(21), I(6) => I6(21), I(7) => I7(21),
    I(8) => I8(21), I(9) => I9(21), I(10) => I10(21), I(11) => I11(21),
    I(12) => I12(21), I(13) => I13(21), I(14) => I14(21), I(15) => I15(21),
    I(16) => I16(21), I(17) => I17(21), I(18) => I18(21), I(19) => I19(21),
    I(20) => I20(21), I(21) => I21(21), I(22) => I22(21), I(23) => I23(21),
    I(24) => I24(21), I(25) => I25(21), I(26) => I26(21), I(27) => I27(21),
    I(28) => I28(21), I(29) => I29(21), I(30) => I30(21), I(31) => I31(21),
    S => S, Y => Y(21));
    
    bit22: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(22), I(1) => I1(22), I(2) => I2(22), I(3) => I3(22),
    I(4) => I4(22), I(5) => I5(22), I(6) => I6(22), I(7) => I7(22),
    I(8) => I8(22), I(9) => I9(22), I(10) => I10(22), I(11) => I11(22),
    I(12) => I12(22), I(13) => I13(22), I(14) => I14(22), I(15) => I15(22),
    I(16) => I16(22), I(17) => I17(22), I(18) => I18(22), I(19) => I19(22),
    I(20) => I20(22), I(21) => I21(22), I(22) => I22(22), I(23) => I23(22),
    I(24) => I24(22), I(25) => I25(22), I(26) => I26(22), I(27) => I27(22),
    I(28) => I28(22), I(29) => I29(22), I(30) => I30(22), I(31) => I31(22),
    S => S, Y => Y(22));
    
    bit23: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(23), I(1) => I1(23), I(2) => I2(23), I(3) => I3(23),
    I(4) => I4(23), I(5) => I5(23), I(6) => I6(23), I(7) => I7(23),
    I(8) => I8(23), I(9) => I9(23), I(10) => I10(23), I(11) => I11(23),
    I(12) => I12(23), I(13) => I13(23), I(14) => I14(23), I(15) => I15(23),
    I(16) => I16(23), I(17) => I17(23), I(18) => I18(23), I(19) => I19(23),
    I(20) => I20(23), I(21) => I21(23), I(22) => I22(23), I(23) => I23(23),
    I(24) => I24(23), I(25) => I25(23), I(26) => I26(23), I(27) => I27(23),
    I(28) => I28(23), I(29) => I29(23), I(30) => I30(23), I(31) => I31(23),
    S => S, Y => Y(23));
    
    bit24: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(24), I(1) => I1(24), I(2) => I2(24), I(3) => I3(24),
    I(4) => I4(24), I(5) => I5(24), I(6) => I6(24), I(7) => I7(24),
    I(8) => I8(24), I(9) => I9(24), I(10) => I10(24), I(11) => I11(24),
    I(12) => I12(24), I(13) => I13(24), I(14) => I14(24), I(15) => I15(24),
    I(16) => I16(24), I(17) => I17(24), I(18) => I18(24), I(19) => I19(24),
    I(20) => I20(24), I(21) => I21(24), I(22) => I22(24), I(23) => I23(24),
    I(24) => I24(24), I(25) => I25(24), I(26) => I26(24), I(27) => I27(24),
    I(28) => I28(24), I(29) => I29(24), I(30) => I30(24), I(31) => I31(24),
    S => S, Y => Y(24));
    
    bit25: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(25), I(1) => I1(25), I(2) => I2(25), I(3) => I3(25),
    I(4) => I4(25), I(5) => I5(25), I(6) => I6(25), I(7) => I7(25),
    I(8) => I8(25), I(9) => I9(25), I(10) => I10(25), I(11) => I11(25),
    I(12) => I12(25), I(13) => I13(25), I(14) => I14(25), I(15) => I15(25),
    I(16) => I16(25), I(17) => I17(25), I(18) => I18(25), I(19) => I19(25),
    I(20) => I20(25), I(21) => I21(25), I(22) => I22(25), I(23) => I23(25),
    I(24) => I24(25), I(25) => I25(25), I(26) => I26(25), I(27) => I27(25),
    I(28) => I28(25), I(29) => I29(25), I(30) => I30(25), I(31) => I31(25),
    S => S, Y => Y(25));
    
    bit26: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(26), I(1) => I1(26), I(2) => I2(26), I(3) => I3(26),
    I(4) => I4(26), I(5) => I5(26), I(6) => I6(26), I(7) => I7(26),
    I(8) => I8(26), I(9) => I9(26), I(10) => I10(26), I(11) => I11(26),
    I(12) => I12(26), I(13) => I13(26), I(14) => I14(26), I(15) => I15(26),
    I(16) => I16(26), I(17) => I17(26), I(18) => I18(26), I(19) => I19(26),
    I(20) => I20(26), I(21) => I21(26), I(22) => I22(26), I(23) => I23(26),
    I(24) => I24(26), I(25) => I25(26), I(26) => I26(26), I(27) => I27(26),
    I(28) => I28(26), I(29) => I29(26), I(30) => I30(26), I(31) => I31(26),
    S => S, Y => Y(26));
    
    bit27: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(27), I(1) => I1(27), I(2) => I2(27), I(3) => I3(27),
    I(4) => I4(27), I(5) => I5(27), I(6) => I6(27), I(7) => I7(27),
    I(8) => I8(27), I(9) => I9(27), I(10) => I10(27), I(11) => I11(27),
    I(12) => I12(27), I(13) => I13(27), I(14) => I14(27), I(15) => I15(27),
    I(16) => I16(27), I(17) => I17(27), I(18) => I18(27), I(19) => I19(27),
    I(20) => I20(27), I(21) => I21(27), I(22) => I22(27), I(23) => I23(27),
    I(24) => I24(27), I(25) => I25(27), I(26) => I26(27), I(27) => I27(27),
    I(28) => I28(27), I(29) => I29(27), I(30) => I30(27), I(31) => I31(27),
    S => S, Y => Y(27));
    
    bit28: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(28), I(1) => I1(28), I(2) => I2(28), I(3) => I3(28),
    I(4) => I4(28), I(5) => I5(28), I(6) => I6(28), I(7) => I7(28),
    I(8) => I8(28), I(9) => I9(28), I(10) => I10(28), I(11) => I11(28),
    I(12) => I12(28), I(13) => I13(28), I(14) => I14(28), I(15) => I15(28),
    I(16) => I16(28), I(17) => I17(28), I(18) => I18(28), I(19) => I19(28),
    I(20) => I20(28), I(21) => I21(28), I(22) => I22(28), I(23) => I23(28),
    I(24) => I24(28), I(25) => I25(28), I(26) => I26(28), I(27) => I27(28),
    I(28) => I28(28), I(29) => I29(28), I(30) => I30(28), I(31) => I31(28),
    S => S, Y => Y(28));
    
    bit29: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(29), I(1) => I1(29), I(2) => I2(29), I(3) => I3(29),
    I(4) => I4(29), I(5) => I5(29), I(6) => I6(29), I(7) => I7(29),
    I(8) => I8(29), I(9) => I9(29), I(10) => I10(29), I(11) => I11(29),
    I(12) => I12(29), I(13) => I13(29), I(14) => I14(29), I(15) => I15(29),
    I(16) => I16(29), I(17) => I17(29), I(18) => I18(29), I(19) => I19(29),
    I(20) => I20(29), I(21) => I21(29), I(22) => I22(29), I(23) => I23(29),
    I(24) => I24(29), I(25) => I25(29), I(26) => I26(29), I(27) => I27(29),
    I(28) => I28(29), I(29) => I29(29), I(30) => I30(29), I(31) => I31(29),
    S => S, Y => Y(29));
    
    bit30: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(30), I(1) => I1(30), I(2) => I2(30), I(3) => I3(30),
    I(4) => I4(30), I(5) => I5(30), I(6) => I6(30), I(7) => I7(30),
    I(8) => I8(30), I(9) => I9(30), I(10) => I10(30), I(11) => I11(30),
    I(12) => I12(30), I(13) => I13(30), I(14) => I14(30), I(15) => I15(30),
    I(16) => I16(30), I(17) => I17(30), I(18) => I18(30), I(19) => I19(30),
    I(20) => I20(30), I(21) => I21(30), I(22) => I22(30), I(23) => I23(30),
    I(24) => I24(30), I(25) => I25(30), I(26) => I26(30), I(27) => I27(30),
    I(28) => I28(30), I(29) => I29(30), I(30) => I30(30), I(31) => I31(30),
    S => S, Y => Y(30));
    
    bit31: RF_Mux32_1Bit_22335824 port map (
    I(0) => I0(31), I(1) => I1(31), I(2) => I2(31), I(3) => I3(31),
    I(4) => I4(31), I(5) => I5(31), I(6) => I6(31), I(7) => I7(31),
    I(8) => I8(31), I(9) => I9(31), I(10) => I10(31), I(11) => I11(31),
    I(12) => I12(31), I(13) => I13(31), I(14) => I14(31), I(15) => I15(31),
    I(16) => I16(31), I(17) => I17(31), I(18) => I18(31), I(19) => I19(31),
    I(20) => I20(31), I(21) => I21(31), I(22) => I22(31), I(23) => I23(31),
    I(24) => I24(31), I(25) => I25(31), I(26) => I26(31), I(27) => I27(31),
    I(28) => I28(31), I(29) => I29(31), I(30) => I30(31), I(31) => I31(31),
    S => S, Y => Y(31));



end Behavioral;
