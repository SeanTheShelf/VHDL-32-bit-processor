----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Sean Conway
-- 
-- Create Date: 20.12.2023 13:00:15
-- Design Name: 
-- Module Name: CPU_RAM_22335824 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;


entity CPU_RAM_22335824 is
    port(
    Clock : in std_logic;
    Address : in std_logic_vector(31 downto 0);
    DataIn : in std_logic_vector(31 downto 0);
    WriteEnable : in std_logic;
    DataOut : out std_logic_vector(31 downto 0)
    );
end CPU_RAM_22335824;

architecture Behavioral of CPU_RAM_22335824 is

type RAM_array is array (0 to 127) of STD_LOGIC_VECTOR (31 downto 0);

signal RAM : RAM_array :=(
X"00000018", -- 0
X"00000019", -- 1
X"0000001A", -- 2
X"0000001B", -- 3
X"0000001C", -- 4
-- 22335824
-- Opcode = digit 3 = 5 
-- DR = digit 2 = 8 
-- SA = digit 1 = 2 
-- SB = digit 0 = 4
--      Opcode            DR      SA      SB
--    "00000000000000101"&"01000"&"00010"&"00101", -- 5
--    "00000000000000110"&"01001"&"00011"&"00110", -- 6
--    "00000000000000111"&"01010"&"00100"&"00111", -- 7
--    "00000000000001000"&"01011"&"00101"&"01000", -- 8
--    "00000000000001001"&"01100"&"00110"&"01001", -- 9
    
X"0000001D", -- 5
X"0000001E", -- 6
X"0000001F", -- 7
X"00000020", -- 8
X"00000021", -- 9 
    
X"00000022", -- 0A
X"00000023", -- 0B
X"00000024", -- 0C
X"00000025", -- 0D
X"00000026", -- 0E
X"00000027", -- 0F
X"00000028", -- 10
X"00000029", -- 11
X"0000002A", -- 12
X"0000002B", -- 13
X"0000002C", -- 14
X"0000002D", -- 15
X"0000002E", -- 16
X"0000002F", -- 17
X"00000030", -- 18
X"00000031", -- 19
X"00000032", -- 1A
X"00000033", -- 1B
X"00000034", -- 1C
X"00000035", -- 1D
X"00000036", -- 1E
X"00000037", -- 1F
X"00000038", -- 20
X"00000039", -- 21
X"0000003A", -- 22
X"0000003B", -- 23
X"0000003C", -- 24
X"0000003D", -- 25
X"0000003E", -- 26
x"0000003F",
X"00000040", -- 27
X"00000041", -- 28
X"00000042", -- 29
X"00000043", -- 2A
X"00000044", -- 2B
X"00000045", -- 2C
X"00000046", -- 2D
X"00000047", -- 2E
X"00000048", -- 2F
X"00000049", -- 30
X"0000004A", -- 31
X"0000004B", -- 32
X"0000004C", -- 33
X"0000004D", -- 34
X"0000004E", -- 35
X"0000004F", -- 36
X"00000050", -- 37
X"00000051", -- 38
X"00000052", -- 39
X"00000053", -- 3A
X"00000054", -- 3B
X"00000055", -- 3C
X"00000056", -- 3D
X"00000057", -- 3E
X"00000058", -- 3F
X"00000059", -- 40
X"0000005A", -- 41
X"0000005B", -- 42
X"0000005C", -- 43
X"0000005D", -- 44
X"0000005E", -- 45
X"0000005F", -- 46
X"00000060", -- 47
X"00000061", -- 48
X"00000062", -- 49
X"00000063", -- 4A
X"00000064", -- 4B
X"00000065", -- 4C
X"00000066", -- 4D
X"00000067", -- 4E
X"00000068", -- 4F
X"00000069", -- 50
X"0000006A", -- 51
X"0000006B", -- 52
X"0000006C", -- 53
X"0000006D", -- 54
X"0000006E", -- 55
X"0000006F", -- 56
X"00000070", -- 57
X"00000071", -- 58
X"00000072", -- 59
X"00000073", -- 5A
X"00000074", -- 5B
X"00000075", -- 5C
X"00000076", -- 5D
X"00000077", -- 5E
X"00000078", -- 5F
X"00000079", -- 60
X"0000007A", -- 61
X"0000007B", -- 62
X"0000007C", -- 63
X"0000007D", -- 64
X"0000007E", -- 65
X"0000007F", -- 66
X"00000080", -- 67
X"00000081", -- 68
X"00000082", -- 69
X"00000083", -- 6A
X"00000084", -- 6B
X"00000085", -- 6C
X"00000086", -- 6D
X"00000087", -- 6E
X"00000088", -- 6F
X"00000089", -- 70
X"0000008A", -- 71
X"0000008B", -- 72
X"0000008C", -- 73
X"0000008D", -- 74
X"0000008E", -- 75
X"0000008F", -- 76
X"00000090", -- 77
X"00000091", -- 78
X"00000092", -- 79
X"00000093", -- 7A
X"00000094", -- 7B
X"00000095", -- 7C
X"00000096", -- 7D
X"00000097" -- 7E
);

begin
process (Clock)
begin
    if Clock'event and Clock='1' then
        if WriteEnable='1' then
            RAM(to_integer(unsigned(Address(6 downto 0)))) <= DataIn after 2ns;
        end if;
     end if;
end process;

DataOut <= RAM(to_integer(unsigned(Address(6 downto 0)))) after 2ns;

end Behavioral;
