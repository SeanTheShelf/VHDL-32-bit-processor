----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Sean Conway
-- 
-- Create Date: 21.12.2023 10:57:58
-- Design Name: 
-- Module Name: CPU_ControlMemory_22335824 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;


entity CPU_ControlMemory_22335824 is
    port ( Address : in std_logic_vector(16 downto 0);
           NA : out std_logic_vector(16 downto 0); -- 34 - 50 
           MS : out std_logic_vector(2 downto 0); -- 31 - 33
           MC : out std_logic; -- 30 
           IL : out std_logic; -- 29 
           PI : out std_logic; -- 28 
           PL : out std_logic; -- 27 
           TD : out std_logic_vector(3 downto 0); -- 23 - 26 
           TA : out std_logic_vector(3 downto 0); -- 19 - 22 
           TB : out std_logic_vector(3 downto 0); -- 15 - 18 
           MB : out std_logic; -- 14 
           FS : out std_logic_vector (4 downto 0); -- 09 - 13 
           MD : out std_logic; -- 08 
           RW : out std_logic; -- 07
           MM : out std_logic; -- 06 
           MW : out std_logic; -- 05 
           RV : out std_logic; -- 04 
           RC : out std_logic; -- 03 
           RN : out std_logic; -- 02 
           RZ : out std_logic; -- 01
           FL : out std_logic  -- 00
           );
end CPU_ControlMemory_22335824;

architecture Behavioral of CPU_ControlMemory_22335824 is

type ROM_array is array(0 to 127) of std_logic_vector(50 downto 0);

signal ROM : ROM_array :=(

    "00000000000000000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'0',
    "00000000000000001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'1',
    "00000000000000010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'0',
    "00000000000000011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'1',
    "00000000000000100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'0',
    "00000000000000101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'1',
    "00000000000000110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'0',
    "00000000000000111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'1',
    "00000000000001000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'0',
    "00000000000001001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'1',
    "00000000000001010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'0',
    "00000000000001011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'1',
    "00000000000001100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'0',
    "00000000000001101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'1',
    "00000000000001110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'0',
    "00000000000001111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'1',
    "00000000000010000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'0',
    "00000000000010001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'1',
    "00000000000010010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'0',
    "00000000000010011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'1',
    "00000000000010100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'0',
    "00000000000010101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'1',
    "00000000000010110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'0',
    "00000000000010111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'1',
    "00000000000011000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'0',
    "00000000000011001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'1',
    "00000000000011010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'0',
    "00000000000011011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'1',
    "00000000000011100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'0',
    "00000000000011101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'1',
    "00000000000011110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'0',
    "00000000000011111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'1',
    "00000000000100000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'0',
    "00000000000100001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'1',
    "00000000000100010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'0',
    "00000000000100011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'1',
    "00000000000100100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'0',
    "00000000000100101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'1',
    "00000000000100110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'0',
    "00000000000100111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'1',
    "00000000000101000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0',
    "00000000000101001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'1',
    "00000000000101010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'0',
    "00000000000101011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'1',
    "00000000000101100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'0',
    "00000000000101101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'1',
    "00000000000101110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'0',
    "00000000000101111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'1',
    "00000000000110000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'0',
    "00000000000110001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'1',
    "00000000000110010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'0',
    "00000000000110011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'1',
    "00000000000110100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'0'&'0',
    "00000000000110101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'0'&'1',
    "00000000000110110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'1'&'0',
    "00000000000110111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'0'&'1'&'1'&'1'&'1',
    "00000000000111000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'0'&'0',
    "00000000000111001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'0'&'1',
    "00000000000111010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'1'&'0',
    "00000000000111011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'0'&'1'&'1',
    "00000000000111100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'0'&'0',
    "00000000000111101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'0'&'1',
    "00000000000111110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'1'&'0',
    "00000000000111111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'0'&'1'&'1'&'1',
    "00000000001000000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'0'&'0',
    "00000000001000001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'0'&'1',
    "00000000001000010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'1'&'0',
    "00000000001000011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'0'&'1'&'1',
    "00000000001000100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'0'&'0',
    "00000000001000101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'0'&'1',
    "00000000001000110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'1'&'0',
    "00000000001000111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'0'&'1'&'1'&'1'&'1'&'1',
    "00000000001001000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'0'&'0',
    "00000000001001001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'0'&'1',
    "00000000001001010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'1'&'0',
    "00000000001001011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'0'&'1'&'1',
    "00000000001001100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'0'&'0',
    "00000000001001101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'0'&'1',
    "00000000001001110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'1'&'0',
    "00000000001001111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'0'&'1'&'1'&'1',
    "00000000001010000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'0'&'0',
    "00000000001010001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'0'&'1',
    "00000000001010010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'1'&'0',
    "00000000001010011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'0'&'1'&'1',
    "00000000001010100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'0'&'0',
    "00000000001010101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'0'&'1',
    "00000000001010110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'1'&'0',
    "00000000001010111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'0'&'1'&'1'&'1'&'1',
    "00000000001011000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'0'&'0',
    "00000000001011001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'0'&'1',
    "00000000001011010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'1'&'0',
    "00000000001011011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'0'&'1'&'1',
    "00000000001011100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'0'&'0',
    "00000000001011101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'0'&'1',
    "00000000001011110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'1'&'0',
    "00000000001011111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'0'&'1'&'1'&'1',
    "00000000001100000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'0'&'0',
    "00000000001100001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'0'&'1',
    "00000000001100010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'1'&'0',
    "00000000001100011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'0'&'1'&'1',
    "00000000001100100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'0'&'0',
    "00000000001100101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'0'&'1',
    "00000000001100110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'1'&'0',
    "00000000001100111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'0'&'1'&'1'&'1'&'1'&'1'&'1'&'1',
    "00000000001101000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&'0',
    "00000000001101001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'0'&'1',
    "00000000001101010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'1'&'0',
    "00000000001101011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'0'&'1'&'1',
    "00000000001101100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'0'&'0',
    "00000000001101101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'0'&'1',
    "00000000001101110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'1'&'0',
    "00000000001101111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'0'&'1'&'1'&'1',
    "00000000001110000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'0'&'0',
    "00000000001110001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'0'&'1',
    "00000000001110010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'1'&'0',
    "00000000001110011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'0'&'1'&'1',
    "00000000001110100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'0'&'0',
    "00000000001110101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'0'&'1',
    "00000000001110110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'1'&'0',
    "00000000001110111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'0'&'1'&'1'&'1'&'1',
    "00000000001111000"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'0'&'0',
    "00000000001111001"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'0'&'1',
    "00000000001111010"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'1'&'0',
    "00000000001111011"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'0'&'1'&'1',
    "00000000001111100"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'0'&'0',
    "00000000001111101"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'0'&'1',
    "00000000001111110"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'1'&'0',
    "00000000001111111"&"000"&'0'&'0'&'0'&'0'&"0000"&"0000"&"0000"&'0'&"00000"&'0'&'1'&'0'&'0'&'1'&'0'&'1'&'1'&'1'
);

signal content_at_address : std_logic_vector(50 downto 0);

begin

content_at_address <= ROM(to_integer(unsigned(Address(6 downto 0)))) after 2ns;

            NA <= content_at_address(50 downto 34);
            MS <= content_at_address(33 downto 31);
            MC <= content_at_address(30);
            IL <= content_at_address(29);
            PI <= content_at_address(28);
            PL <= content_at_address(27);
            TD <= content_at_address(26 downto 23);
            TA <= content_at_address(22 downto 19);
            TB <= content_at_address(18 downto 15);
            MB <= content_at_address(14);
            FS <= content_at_address(13 downto 9);
            MD <= content_at_address(8);
            RW <= content_at_address(7);
            MM <= content_at_address(6);
            MW <= content_at_address(5);
            RV <= content_at_address(4);
            RC <= content_at_address(3);
            RN <= content_at_address(2);
            RZ <= content_at_address(1);
            FL <= content_at_address(0);


end Behavioral;
