----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Sean Conway
-- 
-- Create Date: 22.10.2023 14:47:16
-- Design Name: 
-- Module Name: RF_Mux32_1Bit_22335824_TB - Simulation
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RF_Mux32_1Bit_22335824_TB is
--  Port ( );
end RF_Mux32_1Bit_22335824_TB;

architecture Simulation of RF_Mux32_1Bit_22335824_TB is

    component RF_Mux32_1Bit_22335824
    Port ( I: in std_logic_vector (31 downto 0);
           S: in std_logic_vector (4 downto 0);
           Y: out std_logic
           );
    end component;
    
    signal I_TB : STD_LOGIC_VECTOR (31 downto 0) := (others => '0');
    signal S_TB : STD_LOGIC_VECTOR (4 downto 0) := (others => '0');
    signal Y_TB : std_logic := '0';
    
    constant StudentID : STD_LOGIC_VECTOR (27 downto 0) := x"154D150";

begin

        uut: RF_Mux32_1Bit_22335824 port map (
        I => I_TB,
        S => S_TB,
        Y => Y_TB
        );
        
stim_proc: process
    begin
    
    S_TB <= "00000";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000000001";
    wait for 60ns;
    
    S_TB <= "00001";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000000010";
    wait for 60ns;
    
    S_TB <= "00010";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000000100";
    wait for 60ns;
    
    S_TB <= "00011";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000001000";
    wait for 60ns;
    
    S_TB <= "00100";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000010000";
    wait for 60ns;
    
    S_TB <= "00101";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000000100000";
    wait for 60ns;
    
    S_TB <= "00110";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000001000000";
    wait for 60ns;
    
    S_TB <= "00111";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000010000000";
    wait for 60ns;
    
    S_TB <= "01000";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000000100000000";
    wait for 60ns;
    
    S_TB <= "01001";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000001000000000";
    wait for 60ns;
    
    S_TB <= "01010";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000010000000000";
    wait for 60ns;
    
    S_TB <= "01011";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000000100000000000";
    wait for 60ns;
    
    S_TB <= "01100";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000001000000000000";
    wait for 60ns;
    
    S_TB <= "01101";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000010000000000000";
    wait for 60ns;
    
    S_TB <= "01110";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000000100000000000000";
    wait for 60ns;
    
    S_TB <= "01111";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000001000000000000000";
    wait for 60ns;
    
    S_TB <= "10000";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000010000000000000000";
    wait for 60ns;
    
    S_TB <= "10001";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000000100000000000000000";
    wait for 60ns;
    
    S_TB <= "10010";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000001000000000000000000";
    wait for 60ns;
    
    S_TB <= "10011";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000010000000000000000000";
    wait for 60ns;
    
    S_TB <= "10100";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000000100000000000000000000";
    wait for 60ns;
    
    S_TB <= "10101";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000001000000000000000000000";
    wait for 60ns;
    
    S_TB <= "10110";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000010000000000000000000000";
    wait for 60ns;
    
    S_TB <= "10111";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000000100000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11000";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000001000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11001";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000010000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11010";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00000100000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11011";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00001000000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11100";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00010000000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11101";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "00100000000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11110";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "01000000000000000000000000000000";
    wait for 60ns;
    
    S_TB <= "11111";
    I_TB <= "00000000000000000000000000000000";
    wait for 60ns;
    I_TB <= "10000000000000000000000000000000";
    wait for 60ns;

    end process;


end Simulation;
